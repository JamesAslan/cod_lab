module mul(   
    input  mul_clk,   
    input  resetn,   
    input  mul_signed,
    input [31:0] x,
    input [31:0] y,
    output [63:0] result
    ); 

    wire mul_sign;
    assign mul_sign = mul_signed;
    wire [32:0] A;
    wire [32:0] B;
    assign A = mul_sign ? {x[31],x} : {1'b0,x};
    assign B = mul_sign ? {y[31],y} : {1'b0,y};

    //////////////////////
    //booth
    wire [34:0] B_extend;    //用于booth两位乘法，低位补�?�?0
    assign B_extend = {B[32],B,1'b0};

    wire [63:0] booth_result01;
    wire [63:0] booth_result02;
    wire [63:0] booth_result03;
    wire [63:0] booth_result04;
    wire [63:0] booth_result05;
    wire [63:0] booth_result06;
    wire [63:0] booth_result07;
    wire [63:0] booth_result08;
    wire [63:0] booth_result09;
    wire [63:0] booth_result10;
    wire [63:0] booth_result11;
    wire [63:0] booth_result12;
    wire [63:0] booth_result13;
    wire [63:0] booth_result14;
    wire [63:0] booth_result15;
    wire [63:0] booth_result16;
    wire [63:0] booth_result17;
    
    wire booth_c01;
    wire booth_c02;
    wire booth_c03;
    wire booth_c04;
    wire booth_c05;
    wire booth_c06;
    wire booth_c07;
    wire booth_c08;
    wire booth_c09;
    wire booth_c10;
    wire booth_c11;
    wire booth_c12;
    wire booth_c13;
    wire booth_c14;
    wire booth_c15;
    wire booth_c16;
    wire booth_c17;

    wire [63:0]A_01;
    wire [63:0]A_02;
    wire [63:0]A_03;
    wire [63:0]A_04;
    wire [63:0]A_05;
    wire [63:0]A_06;
    wire [63:0]A_07;
    wire [63:0]A_08;
    wire [63:0]A_09;
    wire [63:0]A_10;
    wire [63:0]A_11;
    wire [63:0]A_12;
    wire [63:0]A_13;
    wire [63:0]A_14;
    wire [63:0]A_15;
    wire [63:0]A_16;
    wire [63:0]A_17;

    assign A_01 = {{31{A[32]}},A};
    assign A_02 = {{29{A[32]}},A,2'b0};  ////?????????????????????
    assign A_03 = {{27{A[32]}},A,4'b0};
    assign A_04 = {{25{A[32]}},A,6'b0};
    assign A_05 = {{23{A[32]}},A,8'b0};
    assign A_06 = {{21{A[32]}},A,10'b0};
    assign A_07 = {{19{A[32]}},A,12'b0};
    assign A_08 = {{17{A[32]}},A,14'b0};
    assign A_09 = {{15{A[32]}},A,16'b0};
    assign A_10 = {{13{A[32]}},A,18'b0};
    assign A_11 = {{11{A[32]}},A,20'b0};
    assign A_12 = {{9{A[32]}},A,22'b0};
    assign A_13 = {{7{A[32]}},A,24'b0};
    assign A_14 = {{5{A[32]}},A,26'b0};
    assign A_15 = {{3{A[32]}},A,28'b0};
    assign A_16 = {{1{A[32]}},A,30'b0};
    assign A_17 = {A,32'b0};

    boothpart booth01(A_01,B_extend[0],B_extend[1],B_extend[2],booth_result01,booth_c01);
    boothpart booth02(A_02,B_extend[2],B_extend[3],B_extend[4],booth_result02,booth_c02);
    boothpart booth03(A_03,B_extend[4],B_extend[5],B_extend[6],booth_result03,booth_c03);
    boothpart booth04(A_04,B_extend[6],B_extend[7],B_extend[8],booth_result04,booth_c04);
    boothpart booth05(A_05,B_extend[8],B_extend[9],B_extend[10],booth_result05,booth_c05);
    boothpart booth06(A_06,B_extend[10],B_extend[11],B_extend[12],booth_result06,booth_c06);
    boothpart booth07(A_07,B_extend[12],B_extend[13],B_extend[14],booth_result07,booth_c07);
    boothpart booth08(A_08,B_extend[14],B_extend[15],B_extend[16],booth_result08,booth_c08);
    boothpart booth09(A_09,B_extend[16],B_extend[17],B_extend[18],booth_result09,booth_c09);
    boothpart booth10(A_10,B_extend[18],B_extend[19],B_extend[20],booth_result10,booth_c10);
    boothpart booth11(A_11,B_extend[20],B_extend[21],B_extend[22],booth_result11,booth_c11);
    boothpart booth12(A_12,B_extend[22],B_extend[23],B_extend[24],booth_result12,booth_c12);
    boothpart booth13(A_13,B_extend[24],B_extend[25],B_extend[26],booth_result13,booth_c13);
    boothpart booth14(A_14,B_extend[26],B_extend[27],B_extend[28],booth_result14,booth_c14);
    boothpart booth15(A_15,B_extend[28],B_extend[29],B_extend[30],booth_result15,booth_c15);
    boothpart booth16(A_16,B_extend[30],B_extend[31],B_extend[32],booth_result16,booth_c16);
    boothpart booth17(A_17,B_extend[32],B_extend[33],B_extend[34],booth_result17,booth_c17);
                         
    ////////////////////////
    //switch
    wire [16:0] w0;
    wire [16:0] w1;
    wire [16:0] w2;
    wire [16:0] w3;
    wire [16:0] w4;
    wire [16:0] w5;
    wire [16:0] w6;
    wire [16:0] w7;
    wire [16:0] w8;
    wire [16:0] w9;
    wire [16:0] w10;
    wire [16:0] w11;
    wire [16:0] w12;
    wire [16:0] w13;
    wire [16:0] w14;
    wire [16:0] w15;
    wire [16:0] w16;
    wire [16:0] w17;
    wire [16:0] w18;
    wire [16:0] w19;
    wire [16:0] w20;
    wire [16:0] w21;
    wire [16:0] w22;
    wire [16:0] w23;
    wire [16:0] w24;
    wire [16:0] w25;
    wire [16:0] w26;
    wire [16:0] w27;
    wire [16:0] w28;
    wire [16:0] w29;
    wire [16:0] w30;
    wire [16:0] w31;
    wire [16:0] w32;
    wire [16:0] w33;
    wire [16:0] w34;
    wire [16:0] w35;
    wire [16:0] w36;
    wire [16:0] w37;
    wire [16:0] w38;
    wire [16:0] w39;
    wire [16:0] w40;
    wire [16:0] w41;
    wire [16:0] w42;
    wire [16:0] w43;
    wire [16:0] w44;
    wire [16:0] w45;
    wire [16:0] w46;
    wire [16:0] w47;
    wire [16:0] w48;
    wire [16:0] w49;
    wire [16:0] w50;
    wire [16:0] w51;
    wire [16:0] w52;
    wire [16:0] w53;
    wire [16:0] w54;
    wire [16:0] w55;
    wire [16:0] w56;
    wire [16:0] w57;
    wire [16:0] w58;
    wire [16:0] w59;
    wire [16:0] w60;
    wire [16:0] w61;
    wire [16:0] w62;
    wire [16:0] w63;


    assign w0 = {booth_result01[0],booth_result02[0],booth_result03[0],booth_result04[0],booth_result05[0],booth_result06[0],booth_result07[0],booth_result08[0],booth_result09[0],booth_result10[0],booth_result11[0],booth_result12[0],booth_result13[0],booth_result14[0],booth_result15[0],booth_result16[0],booth_result17[0]};
    assign w1 = {booth_result01[1],booth_result02[1],booth_result03[1],booth_result04[1],booth_result05[1],booth_result06[1],booth_result07[1],booth_result08[1],booth_result09[1],booth_result10[1],booth_result11[1],booth_result12[1],booth_result13[1],booth_result14[1],booth_result15[1],booth_result16[1],booth_result17[1]};
    assign w2 = {booth_result01[2],booth_result02[2],booth_result03[2],booth_result04[2],booth_result05[2],booth_result06[2],booth_result07[2],booth_result08[2],booth_result09[2],booth_result10[2],booth_result11[2],booth_result12[2],booth_result13[2],booth_result14[2],booth_result15[2],booth_result16[2],booth_result17[2]};
    assign w3 = {booth_result01[3],booth_result02[3],booth_result03[3],booth_result04[3],booth_result05[3],booth_result06[3],booth_result07[3],booth_result08[3],booth_result09[3],booth_result10[3],booth_result11[3],booth_result12[3],booth_result13[3],booth_result14[3],booth_result15[3],booth_result16[3],booth_result17[3]};
    assign w4 = {booth_result01[4],booth_result02[4],booth_result03[4],booth_result04[4],booth_result05[4],booth_result06[4],booth_result07[4],booth_result08[4],booth_result09[4],booth_result10[4],booth_result11[4],booth_result12[4],booth_result13[4],booth_result14[4],booth_result15[4],booth_result16[4],booth_result17[4]};
    assign w5 = {booth_result01[5],booth_result02[5],booth_result03[5],booth_result04[5],booth_result05[5],booth_result06[5],booth_result07[5],booth_result08[5],booth_result09[5],booth_result10[5],booth_result11[5],booth_result12[5],booth_result13[5],booth_result14[5],booth_result15[5],booth_result16[5],booth_result17[5]};
    assign w6 = {booth_result01[6],booth_result02[6],booth_result03[6],booth_result04[6],booth_result05[6],booth_result06[6],booth_result07[6],booth_result08[6],booth_result09[6],booth_result10[6],booth_result11[6],booth_result12[6],booth_result13[6],booth_result14[6],booth_result15[6],booth_result16[6],booth_result17[6]};
    assign w7 = {booth_result01[7],booth_result02[7],booth_result03[7],booth_result04[7],booth_result05[7],booth_result06[7],booth_result07[7],booth_result08[7],booth_result09[7],booth_result10[7],booth_result11[7],booth_result12[7],booth_result13[7],booth_result14[7],booth_result15[7],booth_result16[7],booth_result17[7]};
    assign w8 = {booth_result01[8],booth_result02[8],booth_result03[8],booth_result04[8],booth_result05[8],booth_result06[8],booth_result07[8],booth_result08[8],booth_result09[8],booth_result10[8],booth_result11[8],booth_result12[8],booth_result13[8],booth_result14[8],booth_result15[8],booth_result16[8],booth_result17[8]};
    assign w9 = {booth_result01[9],booth_result02[9],booth_result03[9],booth_result04[9],booth_result05[9],booth_result06[9],booth_result07[9],booth_result08[9],booth_result09[9],booth_result10[9],booth_result11[9],booth_result12[9],booth_result13[9],booth_result14[9],booth_result15[9],booth_result16[9],booth_result17[9]};
    assign w10 = {booth_result01[10],booth_result02[10],booth_result03[10],booth_result04[10],booth_result05[10],booth_result06[10],booth_result07[10],booth_result08[10],booth_result09[10],booth_result10[10],booth_result11[10],booth_result12[10],booth_result13[10],booth_result14[10],booth_result15[10],booth_result16[10],booth_result17[10]};
    assign w11 = {booth_result01[11],booth_result02[11],booth_result03[11],booth_result04[11],booth_result05[11],booth_result06[11],booth_result07[11],booth_result08[11],booth_result09[11],booth_result10[11],booth_result11[11],booth_result12[11],booth_result13[11],booth_result14[11],booth_result15[11],booth_result16[11],booth_result17[11]};
    assign w12 = {booth_result01[12],booth_result02[12],booth_result03[12],booth_result04[12],booth_result05[12],booth_result06[12],booth_result07[12],booth_result08[12],booth_result09[12],booth_result10[12],booth_result11[12],booth_result12[12],booth_result13[12],booth_result14[12],booth_result15[12],booth_result16[12],booth_result17[12]};
    assign w13 = {booth_result01[13],booth_result02[13],booth_result03[13],booth_result04[13],booth_result05[13],booth_result06[13],booth_result07[13],booth_result08[13],booth_result09[13],booth_result10[13],booth_result11[13],booth_result12[13],booth_result13[13],booth_result14[13],booth_result15[13],booth_result16[13],booth_result17[13]};
    assign w14 = {booth_result01[14],booth_result02[14],booth_result03[14],booth_result04[14],booth_result05[14],booth_result06[14],booth_result07[14],booth_result08[14],booth_result09[14],booth_result10[14],booth_result11[14],booth_result12[14],booth_result13[14],booth_result14[14],booth_result15[14],booth_result16[14],booth_result17[14]};
    assign w15 = {booth_result01[15],booth_result02[15],booth_result03[15],booth_result04[15],booth_result05[15],booth_result06[15],booth_result07[15],booth_result08[15],booth_result09[15],booth_result10[15],booth_result11[15],booth_result12[15],booth_result13[15],booth_result14[15],booth_result15[15],booth_result16[15],booth_result17[15]};
    assign w16 = {booth_result01[16],booth_result02[16],booth_result03[16],booth_result04[16],booth_result05[16],booth_result06[16],booth_result07[16],booth_result08[16],booth_result09[16],booth_result10[16],booth_result11[16],booth_result12[16],booth_result13[16],booth_result14[16],booth_result15[16],booth_result16[16],booth_result17[16]};
    assign w17 = {booth_result01[17],booth_result02[17],booth_result03[17],booth_result04[17],booth_result05[17],booth_result06[17],booth_result07[17],booth_result08[17],booth_result09[17],booth_result10[17],booth_result11[17],booth_result12[17],booth_result13[17],booth_result14[17],booth_result15[17],booth_result16[17],booth_result17[17]};
    assign w18 = {booth_result01[18],booth_result02[18],booth_result03[18],booth_result04[18],booth_result05[18],booth_result06[18],booth_result07[18],booth_result08[18],booth_result09[18],booth_result10[18],booth_result11[18],booth_result12[18],booth_result13[18],booth_result14[18],booth_result15[18],booth_result16[18],booth_result17[18]};
    assign w19 = {booth_result01[19],booth_result02[19],booth_result03[19],booth_result04[19],booth_result05[19],booth_result06[19],booth_result07[19],booth_result08[19],booth_result09[19],booth_result10[19],booth_result11[19],booth_result12[19],booth_result13[19],booth_result14[19],booth_result15[19],booth_result16[19],booth_result17[19]};    
    assign w20 = {booth_result01[20],booth_result02[20],booth_result03[20],booth_result04[20],booth_result05[20],booth_result06[20],booth_result07[20],booth_result08[20],booth_result09[20],booth_result10[20],booth_result11[20],booth_result12[20],booth_result13[20],booth_result14[20],booth_result15[20],booth_result16[20],booth_result17[20]};
    assign w21 = {booth_result01[21],booth_result02[21],booth_result03[21],booth_result04[21],booth_result05[21],booth_result06[21],booth_result07[21],booth_result08[21],booth_result09[21],booth_result10[21],booth_result11[21],booth_result12[21],booth_result13[21],booth_result14[21],booth_result15[21],booth_result16[21],booth_result17[21]};
    assign w22 = {booth_result01[22],booth_result02[22],booth_result03[22],booth_result04[22],booth_result05[22],booth_result06[22],booth_result07[22],booth_result08[22],booth_result09[22],booth_result10[22],booth_result11[22],booth_result12[22],booth_result13[22],booth_result14[22],booth_result15[22],booth_result16[22],booth_result17[22]};
    assign w23 = {booth_result01[23],booth_result02[23],booth_result03[23],booth_result04[23],booth_result05[23],booth_result06[23],booth_result07[23],booth_result08[23],booth_result09[23],booth_result10[23],booth_result11[23],booth_result12[23],booth_result13[23],booth_result14[23],booth_result15[23],booth_result16[23],booth_result17[23]};
    assign w24 = {booth_result01[24],booth_result02[24],booth_result03[24],booth_result04[24],booth_result05[24],booth_result06[24],booth_result07[24],booth_result08[24],booth_result09[24],booth_result10[24],booth_result11[24],booth_result12[24],booth_result13[24],booth_result14[24],booth_result15[24],booth_result16[24],booth_result17[24]};
    assign w25 = {booth_result01[25],booth_result02[25],booth_result03[25],booth_result04[25],booth_result05[25],booth_result06[25],booth_result07[25],booth_result08[25],booth_result09[25],booth_result10[25],booth_result11[25],booth_result12[25],booth_result13[25],booth_result14[25],booth_result15[25],booth_result16[25],booth_result17[25]};
    assign w26 = {booth_result01[26],booth_result02[26],booth_result03[26],booth_result04[26],booth_result05[26],booth_result06[26],booth_result07[26],booth_result08[26],booth_result09[26],booth_result10[26],booth_result11[26],booth_result12[26],booth_result13[26],booth_result14[26],booth_result15[26],booth_result16[26],booth_result17[26]};
    assign w27 = {booth_result01[27],booth_result02[27],booth_result03[27],booth_result04[27],booth_result05[27],booth_result06[27],booth_result07[27],booth_result08[27],booth_result09[27],booth_result10[27],booth_result11[27],booth_result12[27],booth_result13[27],booth_result14[27],booth_result15[27],booth_result16[27],booth_result17[27]};
    assign w28 = {booth_result01[28],booth_result02[28],booth_result03[28],booth_result04[28],booth_result05[28],booth_result06[28],booth_result07[28],booth_result08[28],booth_result09[28],booth_result10[28],booth_result11[28],booth_result12[28],booth_result13[28],booth_result14[28],booth_result15[28],booth_result16[28],booth_result17[28]};
    assign w29 = {booth_result01[29],booth_result02[29],booth_result03[29],booth_result04[29],booth_result05[29],booth_result06[29],booth_result07[29],booth_result08[29],booth_result09[29],booth_result10[29],booth_result11[29],booth_result12[29],booth_result13[29],booth_result14[29],booth_result15[29],booth_result16[29],booth_result17[29]};
    assign w30 = {booth_result01[30],booth_result02[30],booth_result03[30],booth_result04[30],booth_result05[30],booth_result06[30],booth_result07[30],booth_result08[30],booth_result09[30],booth_result10[30],booth_result11[30],booth_result12[30],booth_result13[30],booth_result14[30],booth_result15[30],booth_result16[30],booth_result17[30]};
    assign w31 = {booth_result01[31],booth_result02[31],booth_result03[31],booth_result04[31],booth_result05[31],booth_result06[31],booth_result07[31],booth_result08[31],booth_result09[31],booth_result10[31],booth_result11[31],booth_result12[31],booth_result13[31],booth_result14[31],booth_result15[31],booth_result16[31],booth_result17[31]};
    assign w32 = {booth_result01[32],booth_result02[32],booth_result03[32],booth_result04[32],booth_result05[32],booth_result06[32],booth_result07[32],booth_result08[32],booth_result09[32],booth_result10[32],booth_result11[32],booth_result12[32],booth_result13[32],booth_result14[32],booth_result15[32],booth_result16[32],booth_result17[32]};
    assign w33 = {booth_result01[33],booth_result02[33],booth_result03[33],booth_result04[33],booth_result05[33],booth_result06[33],booth_result07[33],booth_result08[33],booth_result09[33],booth_result10[33],booth_result11[33],booth_result12[33],booth_result13[33],booth_result14[33],booth_result15[33],booth_result16[33],booth_result17[33]};
    assign w34 = {booth_result01[34],booth_result02[34],booth_result03[34],booth_result04[34],booth_result05[34],booth_result06[34],booth_result07[34],booth_result08[34],booth_result09[34],booth_result10[34],booth_result11[34],booth_result12[34],booth_result13[34],booth_result14[34],booth_result15[34],booth_result16[34],booth_result17[34]};
    assign w35 = {booth_result01[35],booth_result02[35],booth_result03[35],booth_result04[35],booth_result05[35],booth_result06[35],booth_result07[35],booth_result08[35],booth_result09[35],booth_result10[35],booth_result11[35],booth_result12[35],booth_result13[35],booth_result14[35],booth_result15[35],booth_result16[35],booth_result17[35]};
    assign w36 = {booth_result01[36],booth_result02[36],booth_result03[36],booth_result04[36],booth_result05[36],booth_result06[36],booth_result07[36],booth_result08[36],booth_result09[36],booth_result10[36],booth_result11[36],booth_result12[36],booth_result13[36],booth_result14[36],booth_result15[36],booth_result16[36],booth_result17[36]};
    assign w37 = {booth_result01[37],booth_result02[37],booth_result03[37],booth_result04[37],booth_result05[37],booth_result06[37],booth_result07[37],booth_result08[37],booth_result09[37],booth_result10[37],booth_result11[37],booth_result12[37],booth_result13[37],booth_result14[37],booth_result15[37],booth_result16[37],booth_result17[37]};
    assign w38 = {booth_result01[38],booth_result02[38],booth_result03[38],booth_result04[38],booth_result05[38],booth_result06[38],booth_result07[38],booth_result08[38],booth_result09[38],booth_result10[38],booth_result11[38],booth_result12[38],booth_result13[38],booth_result14[38],booth_result15[38],booth_result16[38],booth_result17[38]};
    assign w39 = {booth_result01[39],booth_result02[39],booth_result03[39],booth_result04[39],booth_result05[39],booth_result06[39],booth_result07[39],booth_result08[39],booth_result09[39],booth_result10[39],booth_result11[39],booth_result12[39],booth_result13[39],booth_result14[39],booth_result15[39],booth_result16[39],booth_result17[39]};
    assign w40 = {booth_result01[40],booth_result02[40],booth_result03[40],booth_result04[40],booth_result05[40],booth_result06[40],booth_result07[40],booth_result08[40],booth_result09[40],booth_result10[40],booth_result11[40],booth_result12[40],booth_result13[40],booth_result14[40],booth_result15[40],booth_result16[40],booth_result17[40]};
    assign w41 = {booth_result01[41],booth_result02[41],booth_result03[41],booth_result04[41],booth_result05[41],booth_result06[41],booth_result07[41],booth_result08[41],booth_result09[41],booth_result10[41],booth_result11[41],booth_result12[41],booth_result13[41],booth_result14[41],booth_result15[41],booth_result16[41],booth_result17[41]};
    assign w42 = {booth_result01[42],booth_result02[42],booth_result03[42],booth_result04[42],booth_result05[42],booth_result06[42],booth_result07[42],booth_result08[42],booth_result09[42],booth_result10[42],booth_result11[42],booth_result12[42],booth_result13[42],booth_result14[42],booth_result15[42],booth_result16[42],booth_result17[42]};
    assign w43 = {booth_result01[43],booth_result02[43],booth_result03[43],booth_result04[43],booth_result05[43],booth_result06[43],booth_result07[43],booth_result08[43],booth_result09[43],booth_result10[43],booth_result11[43],booth_result12[43],booth_result13[43],booth_result14[43],booth_result15[43],booth_result16[43],booth_result17[43]};
    assign w44 = {booth_result01[44],booth_result02[44],booth_result03[44],booth_result04[44],booth_result05[44],booth_result06[44],booth_result07[44],booth_result08[44],booth_result09[44],booth_result10[44],booth_result11[44],booth_result12[44],booth_result13[44],booth_result14[44],booth_result15[44],booth_result16[44],booth_result17[44]};
    assign w45 = {booth_result01[45],booth_result02[45],booth_result03[45],booth_result04[45],booth_result05[45],booth_result06[45],booth_result07[45],booth_result08[45],booth_result09[45],booth_result10[45],booth_result11[45],booth_result12[45],booth_result13[45],booth_result14[45],booth_result15[45],booth_result16[45],booth_result17[45]};
    assign w46 = {booth_result01[46],booth_result02[46],booth_result03[46],booth_result04[46],booth_result05[46],booth_result06[46],booth_result07[46],booth_result08[46],booth_result09[46],booth_result10[46],booth_result11[46],booth_result12[46],booth_result13[46],booth_result14[46],booth_result15[46],booth_result16[46],booth_result17[46]};
    assign w47 = {booth_result01[47],booth_result02[47],booth_result03[47],booth_result04[47],booth_result05[47],booth_result06[47],booth_result07[47],booth_result08[47],booth_result09[47],booth_result10[47],booth_result11[47],booth_result12[47],booth_result13[47],booth_result14[47],booth_result15[47],booth_result16[47],booth_result17[47]};
    assign w48 = {booth_result01[48],booth_result02[48],booth_result03[48],booth_result04[48],booth_result05[48],booth_result06[48],booth_result07[48],booth_result08[48],booth_result09[48],booth_result10[48],booth_result11[48],booth_result12[48],booth_result13[48],booth_result14[48],booth_result15[48],booth_result16[48],booth_result17[48]};
    assign w49 = {booth_result01[49],booth_result02[49],booth_result03[49],booth_result04[49],booth_result05[49],booth_result06[49],booth_result07[49],booth_result08[49],booth_result09[49],booth_result10[49],booth_result11[49],booth_result12[49],booth_result13[49],booth_result14[49],booth_result15[49],booth_result16[49],booth_result17[49]};
    assign w50 = {booth_result01[50],booth_result02[50],booth_result03[50],booth_result04[50],booth_result05[50],booth_result06[50],booth_result07[50],booth_result08[50],booth_result09[50],booth_result10[50],booth_result11[50],booth_result12[50],booth_result13[50],booth_result14[50],booth_result15[50],booth_result16[50],booth_result17[50]};
    assign w51 = {booth_result01[51],booth_result02[51],booth_result03[51],booth_result04[51],booth_result05[51],booth_result06[51],booth_result07[51],booth_result08[51],booth_result09[51],booth_result10[51],booth_result11[51],booth_result12[51],booth_result13[51],booth_result14[51],booth_result15[51],booth_result16[51],booth_result17[51]};
    assign w52 = {booth_result01[52],booth_result02[52],booth_result03[52],booth_result04[52],booth_result05[52],booth_result06[52],booth_result07[52],booth_result08[52],booth_result09[52],booth_result10[52],booth_result11[52],booth_result12[52],booth_result13[52],booth_result14[52],booth_result15[52],booth_result16[52],booth_result17[52]};
    assign w53 = {booth_result01[53],booth_result02[53],booth_result03[53],booth_result04[53],booth_result05[53],booth_result06[53],booth_result07[53],booth_result08[53],booth_result09[53],booth_result10[53],booth_result11[53],booth_result12[53],booth_result13[53],booth_result14[53],booth_result15[53],booth_result16[53],booth_result17[53]};
    assign w54 = {booth_result01[54],booth_result02[54],booth_result03[54],booth_result04[54],booth_result05[54],booth_result06[54],booth_result07[54],booth_result08[54],booth_result09[54],booth_result10[54],booth_result11[54],booth_result12[54],booth_result13[54],booth_result14[54],booth_result15[54],booth_result16[54],booth_result17[54]};
    assign w55 = {booth_result01[55],booth_result02[55],booth_result03[55],booth_result04[55],booth_result05[55],booth_result06[55],booth_result07[55],booth_result08[55],booth_result09[55],booth_result10[55],booth_result11[55],booth_result12[55],booth_result13[55],booth_result14[55],booth_result15[55],booth_result16[55],booth_result17[55]};
    assign w56 = {booth_result01[56],booth_result02[56],booth_result03[56],booth_result04[56],booth_result05[56],booth_result06[56],booth_result07[56],booth_result08[56],booth_result09[56],booth_result10[56],booth_result11[56],booth_result12[56],booth_result13[56],booth_result14[56],booth_result15[56],booth_result16[56],booth_result17[56]};
    assign w57 = {booth_result01[57],booth_result02[57],booth_result03[57],booth_result04[57],booth_result05[57],booth_result06[57],booth_result07[57],booth_result08[57],booth_result09[57],booth_result10[57],booth_result11[57],booth_result12[57],booth_result13[57],booth_result14[57],booth_result15[57],booth_result16[57],booth_result17[57]};
    assign w58 = {booth_result01[58],booth_result02[58],booth_result03[58],booth_result04[58],booth_result05[58],booth_result06[58],booth_result07[58],booth_result08[58],booth_result09[58],booth_result10[58],booth_result11[58],booth_result12[58],booth_result13[58],booth_result14[58],booth_result15[58],booth_result16[58],booth_result17[58]};
    assign w59 = {booth_result01[59],booth_result02[59],booth_result03[59],booth_result04[59],booth_result05[59],booth_result06[59],booth_result07[59],booth_result08[59],booth_result09[59],booth_result10[59],booth_result11[59],booth_result12[59],booth_result13[59],booth_result14[59],booth_result15[59],booth_result16[59],booth_result17[59]};
    assign w60 = {booth_result01[60],booth_result02[60],booth_result03[60],booth_result04[60],booth_result05[60],booth_result06[60],booth_result07[60],booth_result08[60],booth_result09[60],booth_result10[60],booth_result11[60],booth_result12[60],booth_result13[60],booth_result14[60],booth_result15[60],booth_result16[60],booth_result17[60]};
    assign w61 = {booth_result01[61],booth_result02[61],booth_result03[61],booth_result04[61],booth_result05[61],booth_result06[61],booth_result07[61],booth_result08[61],booth_result09[61],booth_result10[61],booth_result11[61],booth_result12[61],booth_result13[61],booth_result14[61],booth_result15[61],booth_result16[61],booth_result17[61]};
    assign w62 = {booth_result01[62],booth_result02[62],booth_result03[62],booth_result04[62],booth_result05[62],booth_result06[62],booth_result07[62],booth_result08[62],booth_result09[62],booth_result10[62],booth_result11[62],booth_result12[62],booth_result13[62],booth_result14[62],booth_result15[62],booth_result16[62],booth_result17[62]};
    assign w63 = {booth_result01[63],booth_result02[63],booth_result03[63],booth_result04[63],booth_result05[63],booth_result06[63],booth_result07[63],booth_result08[63],booth_result09[63],booth_result10[63],booth_result11[63],booth_result12[63],booth_result13[63],booth_result14[63],booth_result15[63],booth_result16[63],booth_result17[63]};

    reg [16:0] w_reg0;
    reg [16:0] w_reg1;
    reg [16:0] w_reg2;
    reg [16:0] w_reg3;
    reg [16:0] w_reg4;
    reg [16:0] w_reg5;
    reg [16:0] w_reg6;
    reg [16:0] w_reg7;
    reg [16:0] w_reg8;
    reg [16:0] w_reg9;
    reg [16:0] w_reg10;
    reg [16:0] w_reg11;
    reg [16:0] w_reg12;
    reg [16:0] w_reg13;
    reg [16:0] w_reg14;
    reg [16:0] w_reg15;
    reg [16:0] w_reg16;
    reg [16:0] w_reg17;
    reg [16:0] w_reg18;
    reg [16:0] w_reg19;
    reg [16:0] w_reg20;
    reg [16:0] w_reg21;
    reg [16:0] w_reg22;
    reg [16:0] w_reg23;
    reg [16:0] w_reg24;
    reg [16:0] w_reg25;
    reg [16:0] w_reg26;
    reg [16:0] w_reg27;
    reg [16:0] w_reg28;
    reg [16:0] w_reg29;
    reg [16:0] w_reg30;
    reg [16:0] w_reg31;
    reg [16:0] w_reg32;
    reg [16:0] w_reg33;
    reg [16:0] w_reg34;
    reg [16:0] w_reg35;
    reg [16:0] w_reg36;
    reg [16:0] w_reg37;
    reg [16:0] w_reg38;
    reg [16:0] w_reg39;
    reg [16:0] w_reg40;
    reg [16:0] w_reg41;
    reg [16:0] w_reg42;
    reg [16:0] w_reg43;
    reg [16:0] w_reg44;
    reg [16:0] w_reg45;
    reg [16:0] w_reg46;
    reg [16:0] w_reg47;
    reg [16:0] w_reg48;
    reg [16:0] w_reg49;
    reg [16:0] w_reg50;
    reg [16:0] w_reg51;
    reg [16:0] w_reg52;
    reg [16:0] w_reg53;
    reg [16:0] w_reg54;
    reg [16:0] w_reg55;
    reg [16:0] w_reg56;
    reg [16:0] w_reg57;
    reg [16:0] w_reg58;
    reg [16:0] w_reg59;
    reg [16:0] w_reg60;
    reg [16:0] w_reg61;
    reg [16:0] w_reg62;
    reg [16:0] w_reg63;

    always @(posedge mul_clk)
	begin
		if(!resetn)
		begin
			w_reg0 <= 17'b0;
            w_reg1 <= 17'b0;
            w_reg2 <= 17'b0;
            w_reg3 <= 17'b0;
            w_reg4 <= 17'b0;
            w_reg5 <= 17'b0;
            w_reg6 <= 17'b0;
            w_reg7 <= 17'b0;
            w_reg8 <= 17'b0;
            w_reg9 <= 17'b0;
            w_reg10 <= 17'b0;
            w_reg11 <= 17'b0;
            w_reg12 <= 17'b0;
            w_reg13 <= 17'b0;
            w_reg14 <= 17'b0;
            w_reg15 <= 17'b0;
            w_reg16 <= 17'b0;
            w_reg17 <= 17'b0;
            w_reg18 <= 17'b0;
            w_reg19 <= 17'b0;
            w_reg20 <= 17'b0;
            w_reg21 <= 17'b0;
            w_reg22 <= 17'b0;
            w_reg23 <= 17'b0;
            w_reg24 <= 17'b0;
            w_reg25 <= 17'b0;
            w_reg26 <= 17'b0;
            w_reg27 <= 17'b0;
            w_reg28 <= 17'b0;
            w_reg29 <= 17'b0;
            w_reg30 <= 17'b0;
            w_reg31 <= 17'b0;
            w_reg32 <= 17'b0;
            w_reg33 <= 17'b0;
            w_reg34 <= 17'b0;
            w_reg35 <= 17'b0;
            w_reg36 <= 17'b0;
            w_reg37 <= 17'b0;
            w_reg38 <= 17'b0;
            w_reg39 <= 17'b0;
            w_reg40 <= 17'b0;
            w_reg41 <= 17'b0;
            w_reg42 <= 17'b0;
            w_reg43 <= 17'b0;
            w_reg44 <= 17'b0;
            w_reg45 <= 17'b0;
            w_reg46 <= 17'b0;
            w_reg47 <= 17'b0;
            w_reg48 <= 17'b0;
            w_reg49 <= 17'b0;
            w_reg50 <= 17'b0;
            w_reg51 <= 17'b0;
            w_reg52 <= 17'b0;
            w_reg53 <= 17'b0;
            w_reg54 <= 17'b0;
            w_reg55 <= 17'b0;
            w_reg56 <= 17'b0;
            w_reg57 <= 17'b0;
            w_reg58 <= 17'b0;
            w_reg59 <= 17'b0;
            w_reg60 <= 17'b0;
            w_reg61 <= 17'b0;
            w_reg62 <= 17'b0;
            w_reg63 <= 17'b0;
            cin0_reg <= 14'b0;
            booth_c15_reg <= 1'b0;
            booth_c16_reg <= 1'b0;
		end
		else
		begin
			w_reg0 <= w0;
            w_reg1 <= w1;
            w_reg2 <= w2;
            w_reg3 <= w3;
            w_reg4 <= w4;
            w_reg5 <= w5;
            w_reg6 <= w6;
            w_reg7 <= w7;
            w_reg8 <= w8;
            w_reg9 <= w9;
            w_reg10 <= w10;
            w_reg11 <= w11;
            w_reg12 <= w12;
            w_reg13 <= w13;
            w_reg14 <= w14;
            w_reg15 <= w15;
            w_reg16 <= w16;
            w_reg17 <= w17;
            w_reg18 <= w18;
            w_reg19 <= w19;
            w_reg20 <= w20;
            w_reg21 <= w21;
            w_reg22 <= w22;
            w_reg23 <= w23;
            w_reg24 <= w24;
            w_reg25 <= w25;
            w_reg26 <= w26;
            w_reg27 <= w27;
            w_reg28 <= w28;
            w_reg29 <= w29;
            w_reg30 <= w30;
            w_reg31 <= w31;
            w_reg32 <= w32;
            w_reg33 <= w33;
            w_reg34 <= w34;
            w_reg35 <= w35;
            w_reg36 <= w36;
            w_reg37 <= w37;
            w_reg38 <= w38;
            w_reg39 <= w39;
            w_reg40 <= w40;
            w_reg41 <= w41;
            w_reg42 <= w42;
            w_reg43 <= w43;
            w_reg44 <= w44;
            w_reg45 <= w45;
            w_reg46 <= w46;
            w_reg47 <= w47;
            w_reg48 <= w48;
            w_reg49 <= w49;
            w_reg50 <= w50;
            w_reg51 <= w51;
            w_reg52 <= w52;
            w_reg53 <= w53;
            w_reg54 <= w54;
            w_reg55 <= w55;
            w_reg56 <= w56;
            w_reg57 <= w57;
            w_reg58 <= w58;
            w_reg59 <= w59;
            w_reg60 <= w60;
            w_reg61 <= w61;
            w_reg62 <= w62;
            w_reg63 <= w63;
            cin0_reg <= cin0;
            booth_c15_reg <= booth_c15;
            booth_c16_reg <= booth_c16;
		end
	end

    reg booth_c16_reg;
    reg booth_c15_reg;
    reg [13:0]cin0_reg;

    ///////////////////////
    //wallace tree
    wire [13:0] cout0;
    wire [13:0] cout1;
    wire [13:0] cout2;
    wire [13:0] cout3;
    wire [13:0] cout4;
    wire [13:0] cout5;
    wire [13:0] cout6;
    wire [13:0] cout7;
    wire [13:0] cout8;
    wire [13:0] cout9;
    wire [13:0] cout10;
    wire [13:0] cout11;
    wire [13:0] cout12;
    wire [13:0] cout13;
    wire [13:0] cout14;
    wire [13:0] cout15;
    wire [13:0] cout16;
    wire [13:0] cout17;
    wire [13:0] cout18;
    wire [13:0] cout19;
    wire [13:0] cout20;
    wire [13:0] cout21;
    wire [13:0] cout22;
    wire [13:0] cout23;
    wire [13:0] cout24;
    wire [13:0] cout25;
    wire [13:0] cout26;
    wire [13:0] cout27;
    wire [13:0] cout28;
    wire [13:0] cout29;
    wire [13:0] cout30;
    wire [13:0] cout31;
    wire [13:0] cout32;
    wire [13:0] cout33;
    wire [13:0] cout34;
    wire [13:0] cout35;
    wire [13:0] cout36;
    wire [13:0] cout37;
    wire [13:0] cout38;
    wire [13:0] cout39;
    wire [13:0] cout40;
    wire [13:0] cout41;
    wire [13:0] cout42;
    wire [13:0] cout43;
    wire [13:0] cout44;
    wire [13:0] cout45;
    wire [13:0] cout46;
    wire [13:0] cout47;
    wire [13:0] cout48;
    wire [13:0] cout49;
    wire [13:0] cout50;
    wire [13:0] cout51;
    wire [13:0] cout52;
    wire [13:0] cout53;
    wire [13:0] cout54;
    wire [13:0] cout55;
    wire [13:0] cout56;
    wire [13:0] cout57;
    wire [13:0] cout58;
    wire [13:0] cout59;
    wire [13:0] cout60;
    wire [13:0] cout61;
    wire [13:0] cout62;
    wire [13:0] cout63;

    wire C0;
    wire C1;
    wire C2;
    wire C3;
    wire C4;
    wire C5;
    wire C6;
    wire C7;
    wire C8;
    wire C9;
    wire C10;
    wire C11;
    wire C12;
    wire C13;
    wire C14;
    wire C15;
    wire C16;
    wire C17;
    wire C18;
    wire C19;
    wire C20;
    wire C21;
    wire C22;
    wire C23;
    wire C24;
    wire C25;
    wire C26;
    wire C27;
    wire C28;
    wire C29;
    wire C30;
    wire C31;
    wire C32;
    wire C33;
    wire C34;
    wire C35;
    wire C36;
    wire C37;
    wire C38;
    wire C39;
    wire C40;
    wire C41;
    wire C42;
    wire C43;
    wire C44;
    wire C45;
    wire C46;
    wire C47;
    wire C48;
    wire C49;
    wire C50;
    wire C51;
    wire C52;
    wire C53;
    wire C54;
    wire C55;
    wire C56;
    wire C57;
    wire C58;
    wire C59;
    wire C60;
    wire C61;
    wire C62;
    wire C63;

    wire S0;
    wire S1;
    wire S2;
    wire S3;
    wire S4;
    wire S5;
    wire S6;
    wire S7;
    wire S8;
    wire S9;
    wire S10;
    wire S11;
    wire S12;
    wire S13;
    wire S14;
    wire S15;
    wire S16;
    wire S17;
    wire S18;
    wire S19;
    wire S20;
    wire S21;
    wire S22;
    wire S23;
    wire S24;
    wire S25;
    wire S26;
    wire S27;
    wire S28;
    wire S29;
    wire S30;
    wire S31;
    wire S32;
    wire S33;
    wire S34;
    wire S35;
    wire S36;
    wire S37;
    wire S38;
    wire S39;
    wire S40;
    wire S41;
    wire S42;
    wire S43;
    wire S44;
    wire S45;
    wire S46;
    wire S47;
    wire S48;
    wire S49;
    wire S50;
    wire S51;
    wire S52;
    wire S53;
    wire S54;
    wire S55;
    wire S56;
    wire S57;
    wire S58;
    wire S59;
    wire S60;
    wire S61;
    wire S62;
    wire S63;

    wire [13:0] cin0;
    assign cin0 = {booth_c01,booth_c02,booth_c03,booth_c04,booth_c05,booth_c06,booth_c07,booth_c08,booth_c09,booth_c10,booth_c11,booth_c12,booth_c13,booth_c14}; 
    
    wallace wallace0(w_reg0,cin0_reg,cout0,C0,S0);
    wallace wallace1(w_reg1,cout0,cout1,C1,S1);
    wallace wallace2(w_reg2,cout1,cout2,C2,S2);
    wallace wallace3(w_reg3,cout2,cout3,C3,S3);
    wallace wallace4(w_reg4,cout3,cout4,C4,S4);
    wallace wallace5(w_reg5,cout4,cout5,C5,S5);
    wallace wallace6(w_reg6,cout5,cout6,C6,S6);
    wallace wallace7(w_reg7,cout6,cout7,C7,S7);
    wallace wallace8(w_reg8,cout7,cout8,C8,S8);
    wallace wallace9(w_reg9,cout8,cout9,C9,S9);
    wallace wallace10(w_reg10,cout9,cout10,C10,S10);
    wallace wallace11(w_reg11,cout10,cout11,C11,S11);
    wallace wallace12(w_reg12,cout11,cout12,C12,S12);
    wallace wallace13(w_reg13,cout12,cout13,C13,S13);
    wallace wallace14(w_reg14,cout13,cout14,C14,S14);
    wallace wallace15(w_reg15,cout14,cout15,C15,S15);
    wallace wallace16(w_reg16,cout15,cout16,C16,S16);
    wallace wallace17(w_reg17,cout16,cout17,C17,S17);
    wallace wallace18(w_reg18,cout17,cout18,C18,S18);
    wallace wallace19(w_reg19,cout18,cout19,C19,S19);
    wallace wallace20(w_reg20,cout19,cout20,C20,S20);
    wallace wallace21(w_reg21,cout20,cout21,C21,S21);
    wallace wallace22(w_reg22,cout21,cout22,C22,S22);
    wallace wallace23(w_reg23,cout22,cout23,C23,S23);
    wallace wallace24(w_reg24,cout23,cout24,C24,S24);
    wallace wallace25(w_reg25,cout24,cout25,C25,S25);
    wallace wallace26(w_reg26,cout25,cout26,C26,S26);
    wallace wallace27(w_reg27,cout26,cout27,C27,S27);
    wallace wallace28(w_reg28,cout27,cout28,C28,S28);
    wallace wallace29(w_reg29,cout28,cout29,C29,S29);
    wallace wallace30(w_reg30,cout29,cout30,C30,S30);
    wallace wallace31(w_reg31,cout30,cout31,C31,S31);
    wallace wallace32(w_reg32,cout31,cout32,C32,S32);
    wallace wallace33(w_reg33,cout32,cout33,C33,S33);
    wallace wallace34(w_reg34,cout33,cout34,C34,S34);
    wallace wallace35(w_reg35,cout34,cout35,C35,S35);
    wallace wallace36(w_reg36,cout35,cout36,C36,S36);
    wallace wallace37(w_reg37,cout36,cout37,C37,S37);
    wallace wallace38(w_reg38,cout37,cout38,C38,S38);
    wallace wallace39(w_reg39,cout38,cout39,C39,S39);
    wallace wallace40(w_reg40,cout39,cout40,C40,S40);
    wallace wallace41(w_reg41,cout40,cout41,C41,S41);
    wallace wallace42(w_reg42,cout41,cout42,C42,S42);
    wallace wallace43(w_reg43,cout42,cout43,C43,S43);
    wallace wallace44(w_reg44,cout43,cout44,C44,S44);
    wallace wallace45(w_reg45,cout44,cout45,C45,S45);
    wallace wallace46(w_reg46,cout45,cout46,C46,S46);
    wallace wallace47(w_reg47,cout46,cout47,C47,S47);
    wallace wallace48(w_reg48,cout47,cout48,C48,S48);
    wallace wallace49(w_reg49,cout48,cout49,C49,S49);
    wallace wallace50(w_reg50,cout49,cout50,C50,S50);
    wallace wallace51(w_reg51,cout50,cout51,C51,S51);
    wallace wallace52(w_reg52,cout51,cout52,C52,S52);
    wallace wallace53(w_reg53,cout52,cout53,C53,S53);
    wallace wallace54(w_reg54,cout53,cout54,C54,S54);
    wallace wallace55(w_reg55,cout54,cout55,C55,S55);
    wallace wallace56(w_reg56,cout55,cout56,C56,S56);
    wallace wallace57(w_reg57,cout56,cout57,C57,S57);
    wallace wallace58(w_reg58,cout57,cout58,C58,S58);
    wallace wallace59(w_reg59,cout58,cout59,C59,S59);
    wallace wallace60(w_reg60,cout59,cout60,C60,S60);
    wallace wallace61(w_reg61,cout60,cout61,C61,S61);
    wallace wallace62(w_reg62,cout61,cout62,C62,S62);
    wallace wallace63(w_reg63,cout62,cout63,C63,S63);

    ////////////////////
    //ADD
    wire [63:0] add_a;
    wire [63:0] add_b;

    assign add_a = {S63,S62,S61,S60,S59,S58,S57,S56,S55,S54,S53,S52,S51,S50,S49,S48,S47,S46,S45,S44,S43,S42,S41,S40,S39,S38,S37,S36,S35,S34,S33,S32,S31,S30,S29,S28,S27,S26,S25,S24,S23,S22,S21,S20,S19,S18,S17,S16,S15,S14,S13,S12,S11,S10,S9,S8,S7,S6,S5,S4,S3,S2,S1,S0};
    assign add_b = {C62,C61,C60,C59,C58,C57,C56,C55,C54,C53,C52,C51,C50,C49,C48,C47,C46,C45,C44,C43,C42,C41,C40,C39,C38,C37,C36,C35,C34,C33,C32,C31,C30,C29,C28,C27,C26,C25,C24,C23,C22,C21,C20,C19,C18,C17,C16,C15,C14,C13,C12,C11,C10,C9,C8,C7,C6,C5,C4,C3,C2,C1,C0,booth_c15_reg};

    assign result = add_a + add_b + booth_c16_reg;

endmodule 
 